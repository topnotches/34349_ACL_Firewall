library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;
entity top_rtl is
  port
  (
    pil_clk : in std_logic;
    pil_rst : in std_logic;

  );
end entity top_rtl;

architecture rtl of top_rtl is

begin

end architecture;