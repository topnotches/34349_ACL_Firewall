library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package ip_packet_pkg is
  type ip_header_rec is record
    ip_header  : std_logic_vector(20 * 4 - 1 downto 0);
    tcp_header : std_logic_vector(20 * 4 - 1 downto 0);
  end record;

  function init_ip_header_rec(
    version          : std_logic_vector(4 - 1 downto 0),
    ihl              : std_logic_vector(4 - 1 downto 0),
    tos              : std_logic_vector(8 - 1 downto 0),
    total_length     : std_logic_vector(16 - 1 downto 0),
    id               : std_logic_vector(16 - 1 downto 0),
    flags_n_frags_os : std_logic_vector(16 - 1 downto 0),
    ttl              : std_logic_vector(8 - 1 downto 0),
    protocol         : std_logic_vector(8 - 1 downto 0),
    head_checksum    : std_logic_vector(16 - 1 downto 0),
    src_addr         : std_logic_vector(32 - 1 downto 0),
    dest_addr        : std_logic_vector(32 - 1 downto 0),
    src_port         : std_logic_vector(16 - 1 downto 0),
    dest_port        : std_logic_vector(16 - 1 downto 0),
    seq_num          : std_logic_vector(32 - 1 downto 0),
    ack_num          : std_logic_vector(32 - 1 downto 0),
    reserved         : std_logic_vector(8 - 1 downto 0),
    flags            : std_logic_vector(8 - 1 downto 0),
    window_size      : std_logic_vector(16 - 1 downto 0),
    checksum         : std_logic_vector(16 - 1 downto 0),
    urgent_pointer   : std_logic_vector(16 - 1 downto 0)
  ) return ip_header_rec;

  function slv_to_ip_header_rec(slv : std_logic_vector) return ip_header_rec;

  function ip_header_rec_to_slv(d_if : ip_header_rec) return std_logic_vector;

end package ip_packet_pkg;

package body ip_packet_pkg is

  function init_ip_header_rec(
    version          : std_logic_vector(4 - 1 downto 0),
    ihl              : std_logic_vector(4 - 1 downto 0),
    tos              : std_logic_vector(8 - 1 downto 0),
    total_length     : std_logic_vector(16 - 1 downto 0),
    id               : std_logic_vector(16 - 1 downto 0),
    flags_n_frags_os : std_logic_vector(16 - 1 downto 0),
    ttl              : std_logic_vector(8 - 1 downto 0),
    protocol         : std_logic_vector(8 - 1 downto 0),
    head_checksum    : std_logic_vector(16 - 1 downto 0),
    src_addr         : std_logic_vector(32 - 1 downto 0),
    dest_addr        : std_logic_vector(32 - 1 downto 0),
    src_port         : std_logic_vector(16 - 1 downto 0),
    dest_port        : std_logic_vector(16 - 1 downto 0),
    seq_num          : std_logic_vector(32 - 1 downto 0),
    ack_num          : std_logic_vector(32 - 1 downto 0),
    reserved         : std_logic_vector(8 - 1 downto 0),
    flags            : std_logic_vector(8 - 1 downto 0),
    window_size      : std_logic_vector(16 - 1 downto 0),
    checksum         : std_logic_vector(16 - 1 downto 0),
    urgent_pointer   : std_logic_vector(16 - 1 downto 0)
  ) return ip_header_rec is
    variable init_data : ip_header_rec;
  begin
    init_data.ip_header  := version & ihl & tos & total_length & id & flags_n_frags_os & ttl & protocol & head_checksum & src_addr & dest_addr;
    init_data.tcp_header := src_port & dest_port & seq_num & ack_num & reserved & flags & window_size & checksum & urgent_pointer;
    return init_data;
  end function init_ip_header_rec;

  function slv_to_ip_header_rec(slv : std_logic_vector) return ip_header_rec is
    variable d_if                     : ip_header_rec;
  begin
    --fill this out
    return d_if
  end slv_to_ip_header_rec;

  function ip_header_rec_to_slv(d_if : ip_header_rec) return std_logic_vector is
    variable slv_result                : std_logic_vector(??);
  begin

    --fill this out
    return slv_result;
  end ip_header_rec_to_slv;

end package body ip_packet_pkg;