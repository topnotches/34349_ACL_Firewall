library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;
use work.acl_defs_pkg.all;

entity hash_table_rtl is
    port
    (
        pil_clk : in std_logic;

        pilv8_hash_table_rd_addr : in std_logic_vector(ACL_HASH_LENGTH - 1 downto 0);
        pil_hash_rd_en           : in std_logic;

        polv128_hash_rd_value : out std_logic_vector(ACL_HASH_TABLE_ADDRESS_LENGTH - 1 downto 0)
        --pilv8_hash_table_wr_addr : in std_logic_vector(ACL_HASH_LENGTH - 1 downto 0);
        --pil_hash_wr_en           : in std_logic;

        --pilv128_hash_wr_value : in std_logic_vector(ACL_HASH_TABLE_ADDRESS_LENGTH - 1 downto 0);
    );
end entity hash_table_rtl;

architecture rtl of hash_table_rtl is
    type hash_table_memory_t is array (0 to ((2 ** ACL_HASH_LENGTH) - 1)) of std_logic_vector(ACL_HASH_TABLE_M9K_LENGTH - 1 downto 0);
    signal sarr256lv32_hash_table_memory_3 : hash_table_memory_t := (-- MSW
    x"00000000", -- 0, 0x00
    x"00000000", -- 1, 0x01
    x"00000000", -- 2, 0x02
    x"00000000", -- 3, 0x03
    x"00000000", -- 4, 0x04
    x"00000000", -- 5, 0x05
    x"00000000", -- 6, 0x06
    x"00000000", -- 7, 0x07
    x"00000000", -- 8, 0x08
    x"00000000", -- 9, 0x09
    x"00000000", -- 10, 0x0a
    x"00000000", -- 11, 0x0b
    x"00000000", -- 12, 0x0c
    x"00000000", -- 13, 0x0d
    x"00000000", -- 14, 0x0e
    x"00000000", -- 15, 0x0f
    x"00000000", -- 16, 0x10
    x"00000000", -- 17, 0x11
    x"00000000", -- 18, 0x12
    x"00000000", -- 19, 0x13
    x"00000000", -- 20, 0x14
    x"00000000", -- 21, 0x15
    x"00000000", -- 22, 0x16
    x"00000000", -- 23, 0x17
    x"00000000", -- 24, 0x18
    x"00000000", -- 25, 0x19
    x"00000000", -- 26, 0x1a
    x"00000000", -- 27, 0x1b
    x"00000000", -- 28, 0x1c
    x"00000000", -- 29, 0x1d
    x"00000000", -- 30, 0x1e
    x"00000000", -- 31, 0x1f
    x"00000000", -- 32, 0x20
    x"00000000", -- 33, 0x21
    x"00000000", -- 34, 0x22
    x"00000000", -- 35, 0x23
    x"00000000", -- 36, 0x24
    x"00000000", -- 37, 0x25
    x"00000000", -- 38, 0x26
    x"00000000", -- 39, 0x27
    x"00000000", -- 40, 0x28
    x"00000000", -- 41, 0x29
    x"00000000", -- 42, 0x2a
    x"00000000", -- 43, 0x2b
    x"00000000", -- 44, 0x2c
    x"00000000", -- 45, 0x2d
    x"00000000", -- 46, 0x2e
    x"00000000", -- 47, 0x2f
    x"00000000", -- 48, 0x30
    x"00000000", -- 49, 0x31
    x"00000000", -- 50, 0x32
    x"00000000", -- 51, 0x33
    x"00000000", -- 52, 0x34
    x"00000000", -- 53, 0x35
    x"00000000", -- 54, 0x36
    x"00000000", -- 55, 0x37
    x"00000000", -- 56, 0x38
    x"00000000", -- 57, 0x39
    x"00000000", -- 58, 0x3a
    x"00000000", -- 59, 0x3b
    x"00000000", -- 60, 0x3c
    x"00000000", -- 61, 0x3d
    x"00000000", -- 62, 0x3e
    x"00000000", -- 63, 0x3f
    x"00000000", -- 64, 0x40
    x"00000000", -- 65, 0x41
    x"00000000", -- 66, 0x42
    x"00000000", -- 67, 0x43
    x"00000000", -- 68, 0x44
    x"00000000", -- 69, 0x45
    x"00000000", -- 70, 0x46
    x"00000000", -- 71, 0x47
    x"00000000", -- 72, 0x48
    x"00000000", -- 73, 0x49
    x"00000000", -- 74, 0x4a
    x"00000000", -- 75, 0x4b
    x"00000000", -- 76, 0x4c
    x"00000000", -- 77, 0x4d
    x"00000000", -- 78, 0x4e
    x"00000000", -- 79, 0x4f
    x"00000000", -- 80, 0x50
    x"00000000", -- 81, 0x51
    x"00000000", -- 82, 0x52
    x"00000000", -- 83, 0x53
    x"00000000", -- 84, 0x54
    x"00000000", -- 85, 0x55
    x"00000000", -- 86, 0x56
    x"00000000", -- 87, 0x57
    x"00000000", -- 88, 0x58
    x"00000000", -- 89, 0x59
    x"00000000", -- 90, 0x5a
    x"00000000", -- 91, 0x5b
    x"00000000", -- 92, 0x5c
    x"00000000", -- 93, 0x5d
    x"00000000", -- 94, 0x5e
    x"00000000", -- 95, 0x5f
    x"00000000", -- 96, 0x60
    x"00000000", -- 97, 0x61
    x"00000000", -- 98, 0x62
    x"00000000", -- 99, 0x63
    x"00000000", -- 100, 0x64
    x"00000000", -- 101, 0x65
    x"00000000", -- 102, 0x66
    x"00000000", -- 103, 0x67
    x"00000000", -- 104, 0x68
    x"00000000", -- 105, 0x69
    x"00000000", -- 106, 0x6a
    x"00000000", -- 107, 0x6b
    x"00000000", -- 108, 0x6c
    x"00000000", -- 109, 0x6d
    x"00000000", -- 110, 0x6e
    x"00000000", -- 111, 0x6f
    x"00000000", -- 112, 0x70
    x"00000000", -- 113, 0x71
    x"00000000", -- 114, 0x72
    x"00000000", -- 115, 0x73
    x"00000000", -- 116, 0x74
    x"00000000", -- 117, 0x75
    x"00000000", -- 118, 0x76
    x"00000000", -- 119, 0x77
    x"00000000", -- 120, 0x78
    x"00000000", -- 121, 0x79
    x"00000000", -- 122, 0x7a
    x"00000000", -- 123, 0x7b
    x"00000000", -- 124, 0x7c
    x"00000000", -- 125, 0x7d
    x"00000000", -- 126, 0x7e
    x"00000000", -- 127, 0x7f
    x"00000000", -- 128, 0x80
    x"00000000", -- 129, 0x81
    x"00000000", -- 130, 0x82
    x"00000000", -- 131, 0x83
    x"00000000", -- 132, 0x84
    x"00000000", -- 133, 0x85
    x"00000000", -- 134, 0x86
    x"00000000", -- 135, 0x87
    x"00000000", -- 136, 0x88
    x"00000000", -- 137, 0x89
    x"00000000", -- 138, 0x8a
    x"00000000", -- 139, 0x8b
    x"00000000", -- 140, 0x8c
    x"00000000", -- 141, 0x8d
    x"00000000", -- 142, 0x8e
    x"00000000", -- 143, 0x8f
    x"00000000", -- 144, 0x90
    x"00000000", -- 145, 0x91
    x"00000000", -- 146, 0x92
    x"00000000", -- 147, 0x93
    x"00000000", -- 148, 0x94
    x"00000000", -- 149, 0x95
    x"00000000", -- 150, 0x96
    x"00000000", -- 151, 0x97
    x"00000000", -- 152, 0x98
    x"00000000", -- 153, 0x99
    x"00000000", -- 154, 0x9a
    x"00000000", -- 155, 0x9b
    x"00000000", -- 156, 0x9c
    x"00000000", -- 157, 0x9d
    x"00000000", -- 158, 0x9e
    x"00000000", -- 159, 0x9f
    x"00000000", -- 160, 0xa0
    x"00000000", -- 161, 0xa1
    x"00000000", -- 162, 0xa2
    x"00000000", -- 163, 0xa3
    x"00000000", -- 164, 0xa4
    x"00000000", -- 165, 0xa5
    x"00000000", -- 166, 0xa6
    x"00000000", -- 167, 0xa7
    x"00000000", -- 168, 0xa8
    x"00000000", -- 169, 0xa9
    x"00000000", -- 170, 0xaa
    x"00000000", -- 171, 0xab
    x"00000000", -- 172, 0xac
    x"00000000", -- 173, 0xad
    x"00000000", -- 174, 0xae
    x"00000000", -- 175, 0xaf
    x"00000000", -- 176, 0xb0
    x"00000000", -- 177, 0xb1
    x"00000000", -- 178, 0xb2
    x"00000000", -- 179, 0xb3
    x"00000000", -- 180, 0xb4
    x"00000000", -- 181, 0xb5
    x"00000000", -- 182, 0xb6
    x"00000000", -- 183, 0xb7
    x"00000000", -- 184, 0xb8
    x"00000000", -- 185, 0xb9
    x"00000000", -- 186, 0xba
    x"00000000", -- 187, 0xbb
    x"00000000", -- 188, 0xbc
    x"00000000", -- 189, 0xbd
    x"00000000", -- 190, 0xbe
    x"00000000", -- 191, 0xbf
    x"00000000", -- 192, 0xc0
    x"00000000", -- 193, 0xc1
    x"00000000", -- 194, 0xc2
    x"00000000", -- 195, 0xc3
    x"00000000", -- 196, 0xc4
    x"00000000", -- 197, 0xc5
    x"00000000", -- 198, 0xc6
    x"F2012345", -- 199, 0xc7
    x"00000000", -- 200, 0xc8
    x"00000000", -- 201, 0xc9
    x"00000000", -- 202, 0xca
    x"00000000", -- 203, 0xcb
    x"00000000", -- 204, 0xcc
    x"00000000", -- 205, 0xcd
    x"00000000", -- 206, 0xce
    x"00000000", -- 207, 0xcf
    x"00000000", -- 208, 0xd0
    x"00000000", -- 209, 0xd1
    x"00000000", -- 210, 0xd2
    x"00000000", -- 211, 0xd3
    x"00000000", -- 212, 0xd4
    x"00000000", -- 213, 0xd5
    x"00000000", -- 214, 0xd6
    x"00000000", -- 215, 0xd7
    x"00000000", -- 216, 0xd8
    x"00000000", -- 217, 0xd9
    x"00000000", -- 218, 0xda
    x"00000000", -- 219, 0xdb
    x"00000000", -- 220, 0xdc
    x"00000000", -- 221, 0xdd
    x"00000000", -- 222, 0xde
    x"00000000", -- 223, 0xdf
    x"00000000", -- 224, 0xe0
    x"00000000", -- 225, 0xe1
    x"3FFFFFFF", -- 226, 0xe2
    x"00000000", -- 227, 0xe3
    x"00000000", -- 228, 0xe4
    x"00000000", -- 229, 0xe5
    x"00000000", -- 230, 0xe6
    x"00000000", -- 231, 0xe7
    x"00000000", -- 232, 0xe8
    x"00000000", -- 233, 0xe9
    x"00000000", -- 234, 0xea
    x"00000000", -- 235, 0xeb
    x"00000000", -- 236, 0xec
    x"00000000", -- 237, 0xed
    x"00000000", -- 238, 0xee
    x"00000000", -- 239, 0xef
    x"00000000", -- 240, 0xf0
    x"00000000", -- 241, 0xf1
    x"00000000", -- 242, 0xf2
    x"00000000", -- 243, 0xf3
    x"00000000", -- 244, 0xf4
    x"00000000", -- 245, 0xf5
    x"00000000", -- 246, 0xf6
    x"00000000", -- 247, 0xf7
    x"00000000", -- 248, 0xf8
    x"00000000", -- 249, 0xf9
    x"00000000", -- 250, 0xfa
    x"00000000", -- 251, 0xfb
    x"00000000", -- 252, 0xfc
    x"00000000", -- 253, 0xfd
    x"00000000", -- 254, 0xfe
    x"00000000" -- 255, 0xff
    );
    signal sarr256lv32_hash_table_memory_2 : hash_table_memory_t := (-- AMSW
    x"00000000", -- 0, 0x00
    x"00000000", -- 1, 0x01
    x"00000000", -- 2, 0x02
    x"00000000", -- 3, 0x03
    x"00000000", -- 4, 0x04
    x"00000000", -- 5, 0x05
    x"00000000", -- 6, 0x06
    x"00000000", -- 7, 0x07
    x"00000000", -- 8, 0x08
    x"00000000", -- 9, 0x09
    x"00000000", -- 10, 0x0a
    x"00000000", -- 11, 0x0b
    x"00000000", -- 12, 0x0c
    x"00000000", -- 13, 0x0d
    x"00000000", -- 14, 0x0e
    x"00000000", -- 15, 0x0f
    x"00000000", -- 16, 0x10
    x"00000000", -- 17, 0x11
    x"00000000", -- 18, 0x12
    x"00000000", -- 19, 0x13
    x"00000000", -- 20, 0x14
    x"00000000", -- 21, 0x15
    x"00000000", -- 22, 0x16
    x"00000000", -- 23, 0x17
    x"00000000", -- 24, 0x18
    x"00000000", -- 25, 0x19
    x"00000000", -- 26, 0x1a
    x"00000000", -- 27, 0x1b
    x"00000000", -- 28, 0x1c
    x"00000000", -- 29, 0x1d
    x"00000000", -- 30, 0x1e
    x"00000000", -- 31, 0x1f
    x"00000000", -- 32, 0x20
    x"00000000", -- 33, 0x21
    x"00000000", -- 34, 0x22
    x"00000000", -- 35, 0x23
    x"00000000", -- 36, 0x24
    x"00000000", -- 37, 0x25
    x"00000000", -- 38, 0x26
    x"00000000", -- 39, 0x27
    x"00000000", -- 40, 0x28
    x"00000000", -- 41, 0x29
    x"00000000", -- 42, 0x2a
    x"00000000", -- 43, 0x2b
    x"00000000", -- 44, 0x2c
    x"00000000", -- 45, 0x2d
    x"00000000", -- 46, 0x2e
    x"00000000", -- 47, 0x2f
    x"00000000", -- 48, 0x30
    x"00000000", -- 49, 0x31
    x"00000000", -- 50, 0x32
    x"00000000", -- 51, 0x33
    x"00000000", -- 52, 0x34
    x"00000000", -- 53, 0x35
    x"00000000", -- 54, 0x36
    x"00000000", -- 55, 0x37
    x"00000000", -- 56, 0x38
    x"00000000", -- 57, 0x39
    x"00000000", -- 58, 0x3a
    x"00000000", -- 59, 0x3b
    x"00000000", -- 60, 0x3c
    x"00000000", -- 61, 0x3d
    x"00000000", -- 62, 0x3e
    x"00000000", -- 63, 0x3f
    x"00000000", -- 64, 0x40
    x"00000000", -- 65, 0x41
    x"00000000", -- 66, 0x42
    x"00000000", -- 67, 0x43
    x"00000000", -- 68, 0x44
    x"00000000", -- 69, 0x45
    x"00000000", -- 70, 0x46
    x"00000000", -- 71, 0x47
    x"00000000", -- 72, 0x48
    x"00000000", -- 73, 0x49
    x"00000000", -- 74, 0x4a
    x"00000000", -- 75, 0x4b
    x"00000000", -- 76, 0x4c
    x"00000000", -- 77, 0x4d
    x"00000000", -- 78, 0x4e
    x"00000000", -- 79, 0x4f
    x"00000000", -- 80, 0x50
    x"00000000", -- 81, 0x51
    x"00000000", -- 82, 0x52
    x"00000000", -- 83, 0x53
    x"00000000", -- 84, 0x54
    x"00000000", -- 85, 0x55
    x"00000000", -- 86, 0x56
    x"00000000", -- 87, 0x57
    x"00000000", -- 88, 0x58
    x"00000000", -- 89, 0x59
    x"00000000", -- 90, 0x5a
    x"00000000", -- 91, 0x5b
    x"00000000", -- 92, 0x5c
    x"00000000", -- 93, 0x5d
    x"00000000", -- 94, 0x5e
    x"00000000", -- 95, 0x5f
    x"00000000", -- 96, 0x60
    x"00000000", -- 97, 0x61
    x"00000000", -- 98, 0x62
    x"00000000", -- 99, 0x63
    x"00000000", -- 100, 0x64
    x"00000000", -- 101, 0x65
    x"00000000", -- 102, 0x66
    x"00000000", -- 103, 0x67
    x"00000000", -- 104, 0x68
    x"00000000", -- 105, 0x69
    x"00000000", -- 106, 0x6a
    x"00000000", -- 107, 0x6b
    x"00000000", -- 108, 0x6c
    x"00000000", -- 109, 0x6d
    x"00000000", -- 110, 0x6e
    x"00000000", -- 111, 0x6f
    x"00000000", -- 112, 0x70
    x"00000000", -- 113, 0x71
    x"00000000", -- 114, 0x72
    x"00000000", -- 115, 0x73
    x"00000000", -- 116, 0x74
    x"00000000", -- 117, 0x75
    x"00000000", -- 118, 0x76
    x"00000000", -- 119, 0x77
    x"00000000", -- 120, 0x78
    x"00000000", -- 121, 0x79
    x"00000000", -- 122, 0x7a
    x"00000000", -- 123, 0x7b
    x"00000000", -- 124, 0x7c
    x"00000000", -- 125, 0x7d
    x"00000000", -- 126, 0x7e
    x"00000000", -- 127, 0x7f
    x"00000000", -- 128, 0x80
    x"00000000", -- 129, 0x81
    x"00000000", -- 130, 0x82
    x"00000000", -- 131, 0x83
    x"00000000", -- 132, 0x84
    x"00000000", -- 133, 0x85
    x"00000000", -- 134, 0x86
    x"00000000", -- 135, 0x87
    x"00000000", -- 136, 0x88
    x"00000000", -- 137, 0x89
    x"00000000", -- 138, 0x8a
    x"00000000", -- 139, 0x8b
    x"00000000", -- 140, 0x8c
    x"00000000", -- 141, 0x8d
    x"00000000", -- 142, 0x8e
    x"00000000", -- 143, 0x8f
    x"00000000", -- 144, 0x90
    x"00000000", -- 145, 0x91
    x"00000000", -- 146, 0x92
    x"00000000", -- 147, 0x93
    x"00000000", -- 148, 0x94
    x"00000000", -- 149, 0x95
    x"00000000", -- 150, 0x96
    x"00000000", -- 151, 0x97
    x"00000000", -- 152, 0x98
    x"00000000", -- 153, 0x99
    x"00000000", -- 154, 0x9a
    x"00000000", -- 155, 0x9b
    x"00000000", -- 156, 0x9c
    x"00000000", -- 157, 0x9d
    x"00000000", -- 158, 0x9e
    x"00000000", -- 159, 0x9f
    x"00000000", -- 160, 0xa0
    x"00000000", -- 161, 0xa1
    x"00000000", -- 162, 0xa2
    x"00000000", -- 163, 0xa3
    x"00000000", -- 164, 0xa4
    x"00000000", -- 165, 0xa5
    x"00000000", -- 166, 0xa6
    x"00000000", -- 167, 0xa7
    x"00000000", -- 168, 0xa8
    x"00000000", -- 169, 0xa9
    x"00000000", -- 170, 0xaa
    x"00000000", -- 171, 0xab
    x"00000000", -- 172, 0xac
    x"00000000", -- 173, 0xad
    x"00000000", -- 174, 0xae
    x"00000000", -- 175, 0xaf
    x"00000000", -- 176, 0xb0
    x"00000000", -- 177, 0xb1
    x"00000000", -- 178, 0xb2
    x"00000000", -- 179, 0xb3
    x"00000000", -- 180, 0xb4
    x"00000000", -- 181, 0xb5
    x"00000000", -- 182, 0xb6
    x"00000000", -- 183, 0xb7
    x"00000000", -- 184, 0xb8
    x"00000000", -- 185, 0xb9
    x"00000000", -- 186, 0xba
    x"00000000", -- 187, 0xbb
    x"00000000", -- 188, 0xbc
    x"00000000", -- 189, 0xbd
    x"00000000", -- 190, 0xbe
    x"00000000", -- 191, 0xbf
    x"00000000", -- 192, 0xc0
    x"00000000", -- 193, 0xc1
    x"00000000", -- 194, 0xc2
    x"00000000", -- 195, 0xc3
    x"00000000", -- 196, 0xc4
    x"00000000", -- 197, 0xc5
    x"00000000", -- 198, 0xc6
    x"6789ABCD", -- 199, 0xc7
    x"00000000", -- 200, 0xc8
    x"00000000", -- 201, 0xc9
    x"00000000", -- 202, 0xca
    x"00000000", -- 203, 0xcb
    x"00000000", -- 204, 0xcc
    x"00000000", -- 205, 0xcd
    x"00000000", -- 206, 0xce
    x"00000000", -- 207, 0xcf
    x"00000000", -- 208, 0xd0
    x"00000000", -- 209, 0xd1
    x"00000000", -- 210, 0xd2
    x"00000000", -- 211, 0xd3
    x"00000000", -- 212, 0xd4
    x"00000000", -- 213, 0xd5
    x"00000000", -- 214, 0xd6
    x"00000000", -- 215, 0xd7
    x"00000000", -- 216, 0xd8
    x"00000000", -- 217, 0xd9
    x"00000000", -- 218, 0xda
    x"00000000", -- 219, 0xdb
    x"00000000", -- 220, 0xdc
    x"00000000", -- 221, 0xdd
    x"00000000", -- 222, 0xde
    x"00000000", -- 223, 0xdf
    x"00000000", -- 224, 0xe0
    x"00000000", -- 225, 0xe1
    x"FFF1FFF1", -- 226, 0xe2
    x"00000000", -- 227, 0xe3
    x"00000000", -- 228, 0xe4
    x"00000000", -- 229, 0xe5
    x"00000000", -- 230, 0xe6
    x"00000000", -- 231, 0xe7
    x"00000000", -- 232, 0xe8
    x"00000000", -- 233, 0xe9
    x"00000000", -- 234, 0xea
    x"00000000", -- 235, 0xeb
    x"00000000", -- 236, 0xec
    x"00000000", -- 237, 0xed
    x"00000000", -- 238, 0xee
    x"00000000", -- 239, 0xef
    x"00000000", -- 240, 0xf0
    x"00000000", -- 241, 0xf1
    x"00000000", -- 242, 0xf2
    x"00000000", -- 243, 0xf3
    x"00000000", -- 244, 0xf4
    x"00000000", -- 245, 0xf5
    x"00000000", -- 246, 0xf6
    x"00000000", -- 247, 0xf7
    x"00000000", -- 248, 0xf8
    x"00000000", -- 249, 0xf9
    x"00000000", -- 250, 0xfa
    x"00000000", -- 251, 0xfb
    x"00000000", -- 252, 0xfc
    x"00000000", -- 253, 0xfd
    x"00000000", -- 254, 0xfe
    x"00000000" -- 255, 0xff

    );
    signal sarr256lv32_hash_table_memory_1 : hash_table_memory_t := (-- ALSW
    x"00000000", -- 0, 0x00
    x"00000000", -- 1, 0x01
    x"00000000", -- 2, 0x02
    x"00000000", -- 3, 0x03
    x"00000000", -- 4, 0x04
    x"00000000", -- 5, 0x05
    x"00000000", -- 6, 0x06
    x"00000000", -- 7, 0x07
    x"00000000", -- 8, 0x08
    x"00000000", -- 9, 0x09
    x"00000000", -- 10, 0x0a
    x"00000000", -- 11, 0x0b
    x"00000000", -- 12, 0x0c
    x"00000000", -- 13, 0x0d
    x"00000000", -- 14, 0x0e
    x"00000000", -- 15, 0x0f
    x"00000000", -- 16, 0x10
    x"00000000", -- 17, 0x11
    x"00000000", -- 18, 0x12
    x"00000000", -- 19, 0x13
    x"00000000", -- 20, 0x14
    x"00000000", -- 21, 0x15
    x"00000000", -- 22, 0x16
    x"00000000", -- 23, 0x17
    x"00000000", -- 24, 0x18
    x"00000000", -- 25, 0x19
    x"00000000", -- 26, 0x1a
    x"00000000", -- 27, 0x1b
    x"00000000", -- 28, 0x1c
    x"00000000", -- 29, 0x1d
    x"00000000", -- 30, 0x1e
    x"00000000", -- 31, 0x1f
    x"00000000", -- 32, 0x20
    x"00000000", -- 33, 0x21
    x"00000000", -- 34, 0x22
    x"00000000", -- 35, 0x23
    x"00000000", -- 36, 0x24
    x"00000000", -- 37, 0x25
    x"00000000", -- 38, 0x26
    x"00000000", -- 39, 0x27
    x"00000000", -- 40, 0x28
    x"00000000", -- 41, 0x29
    x"00000000", -- 42, 0x2a
    x"00000000", -- 43, 0x2b
    x"00000000", -- 44, 0x2c
    x"00000000", -- 45, 0x2d
    x"00000000", -- 46, 0x2e
    x"00000000", -- 47, 0x2f
    x"00000000", -- 48, 0x30
    x"00000000", -- 49, 0x31
    x"00000000", -- 50, 0x32
    x"00000000", -- 51, 0x33
    x"00000000", -- 52, 0x34
    x"00000000", -- 53, 0x35
    x"00000000", -- 54, 0x36
    x"00000000", -- 55, 0x37
    x"00000000", -- 56, 0x38
    x"00000000", -- 57, 0x39
    x"00000000", -- 58, 0x3a
    x"00000000", -- 59, 0x3b
    x"00000000", -- 60, 0x3c
    x"00000000", -- 61, 0x3d
    x"00000000", -- 62, 0x3e
    x"00000000", -- 63, 0x3f
    x"00000000", -- 64, 0x40
    x"00000000", -- 65, 0x41
    x"00000000", -- 66, 0x42
    x"00000000", -- 67, 0x43
    x"00000000", -- 68, 0x44
    x"00000000", -- 69, 0x45
    x"00000000", -- 70, 0x46
    x"00000000", -- 71, 0x47
    x"00000000", -- 72, 0x48
    x"00000000", -- 73, 0x49
    x"00000000", -- 74, 0x4a
    x"00000000", -- 75, 0x4b
    x"00000000", -- 76, 0x4c
    x"00000000", -- 77, 0x4d
    x"00000000", -- 78, 0x4e
    x"00000000", -- 79, 0x4f
    x"00000000", -- 80, 0x50
    x"00000000", -- 81, 0x51
    x"00000000", -- 82, 0x52
    x"00000000", -- 83, 0x53
    x"00000000", -- 84, 0x54
    x"00000000", -- 85, 0x55
    x"00000000", -- 86, 0x56
    x"00000000", -- 87, 0x57
    x"00000000", -- 88, 0x58
    x"00000000", -- 89, 0x59
    x"00000000", -- 90, 0x5a
    x"00000000", -- 91, 0x5b
    x"00000000", -- 92, 0x5c
    x"00000000", -- 93, 0x5d
    x"00000000", -- 94, 0x5e
    x"00000000", -- 95, 0x5f
    x"00000000", -- 96, 0x60
    x"00000000", -- 97, 0x61
    x"00000000", -- 98, 0x62
    x"00000000", -- 99, 0x63
    x"00000000", -- 100, 0x64
    x"00000000", -- 101, 0x65
    x"00000000", -- 102, 0x66
    x"00000000", -- 103, 0x67
    x"00000000", -- 104, 0x68
    x"00000000", -- 105, 0x69
    x"00000000", -- 106, 0x6a
    x"00000000", -- 107, 0x6b
    x"00000000", -- 108, 0x6c
    x"00000000", -- 109, 0x6d
    x"00000000", -- 110, 0x6e
    x"00000000", -- 111, 0x6f
    x"00000000", -- 112, 0x70
    x"00000000", -- 113, 0x71
    x"00000000", -- 114, 0x72
    x"00000000", -- 115, 0x73
    x"00000000", -- 116, 0x74
    x"00000000", -- 117, 0x75
    x"00000000", -- 118, 0x76
    x"00000000", -- 119, 0x77
    x"00000000", -- 120, 0x78
    x"00000000", -- 121, 0x79
    x"00000000", -- 122, 0x7a
    x"00000000", -- 123, 0x7b
    x"00000000", -- 124, 0x7c
    x"00000000", -- 125, 0x7d
    x"00000000", -- 126, 0x7e
    x"00000000", -- 127, 0x7f
    x"00000000", -- 128, 0x80
    x"00000000", -- 129, 0x81
    x"00000000", -- 130, 0x82
    x"00000000", -- 131, 0x83
    x"00000000", -- 132, 0x84
    x"00000000", -- 133, 0x85
    x"00000000", -- 134, 0x86
    x"00000000", -- 135, 0x87
    x"00000000", -- 136, 0x88
    x"00000000", -- 137, 0x89
    x"00000000", -- 138, 0x8a
    x"00000000", -- 139, 0x8b
    x"00000000", -- 140, 0x8c
    x"00000000", -- 141, 0x8d
    x"00000000", -- 142, 0x8e
    x"00000000", -- 143, 0x8f
    x"00000000", -- 144, 0x90
    x"00000000", -- 145, 0x91
    x"00000000", -- 146, 0x92
    x"00000000", -- 147, 0x93
    x"00000000", -- 148, 0x94
    x"00000000", -- 149, 0x95
    x"00000000", -- 150, 0x96
    x"00000000", -- 151, 0x97
    x"00000000", -- 152, 0x98
    x"00000000", -- 153, 0x99
    x"00000000", -- 154, 0x9a
    x"00000000", -- 155, 0x9b
    x"00000000", -- 156, 0x9c
    x"00000000", -- 157, 0x9d
    x"00000000", -- 158, 0x9e
    x"00000000", -- 159, 0x9f
    x"00000000", -- 160, 0xa0
    x"00000000", -- 161, 0xa1
    x"00000000", -- 162, 0xa2
    x"00000000", -- 163, 0xa3
    x"00000000", -- 164, 0xa4
    x"00000000", -- 165, 0xa5
    x"00000000", -- 166, 0xa6
    x"00000000", -- 167, 0xa7
    x"00000000", -- 168, 0xa8
    x"00000000", -- 169, 0xa9
    x"00000000", -- 170, 0xaa
    x"00000000", -- 171, 0xab
    x"00000000", -- 172, 0xac
    x"00000000", -- 173, 0xad
    x"00000000", -- 174, 0xae
    x"00000000", -- 175, 0xaf
    x"00000000", -- 176, 0xb0
    x"00000000", -- 177, 0xb1
    x"00000000", -- 178, 0xb2
    x"00000000", -- 179, 0xb3
    x"00000000", -- 180, 0xb4
    x"00000000", -- 181, 0xb5
    x"00000000", -- 182, 0xb6
    x"00000000", -- 183, 0xb7
    x"00000000", -- 184, 0xb8
    x"00000000", -- 185, 0xb9
    x"00000000", -- 186, 0xba
    x"00000000", -- 187, 0xbb
    x"00000000", -- 188, 0xbc
    x"00000000", -- 189, 0xbd
    x"00000000", -- 190, 0xbe
    x"00000000", -- 191, 0xbf
    x"00000000", -- 192, 0xc0
    x"00000000", -- 193, 0xc1
    x"00000000", -- 194, 0xc2
    x"00000000", -- 195, 0xc3
    x"00000000", -- 196, 0xc4
    x"00000000", -- 197, 0xc5
    x"00000000", -- 198, 0xc6
    x"EF012345", -- 199, 0xc7
    x"00000000", -- 200, 0xc8
    x"00000000", -- 201, 0xc9
    x"00000000", -- 202, 0xca
    x"00000000", -- 203, 0xcb
    x"00000000", -- 204, 0xcc
    x"00000000", -- 205, 0xcd
    x"00000000", -- 206, 0xce
    x"00000000", -- 207, 0xcf
    x"00000000", -- 208, 0xd0
    x"00000000", -- 209, 0xd1
    x"00000000", -- 210, 0xd2
    x"00000000", -- 211, 0xd3
    x"00000000", -- 212, 0xd4
    x"00000000", -- 213, 0xd5
    x"00000000", -- 214, 0xd6
    x"00000000", -- 215, 0xd7
    x"00000000", -- 216, 0xd8
    x"00000000", -- 217, 0xd9
    x"00000000", -- 218, 0xda
    x"00000000", -- 219, 0xdb
    x"00000000", -- 220, 0xdc
    x"00000000", -- 221, 0xdd
    x"00000000", -- 222, 0xde
    x"00000000", -- 223, 0xdf
    x"00000000", -- 224, 0xe0
    x"00000000", -- 225, 0xe1
    x"FFFFFFFF", -- 226, 0xe2
    x"00000000", -- 227, 0xe3
    x"00000000", -- 228, 0xe4
    x"00000000", -- 229, 0xe5
    x"00000000", -- 230, 0xe6
    x"00000000", -- 231, 0xe7
    x"00000000", -- 232, 0xe8
    x"00000000", -- 233, 0xe9
    x"00000000", -- 234, 0xea
    x"00000000", -- 235, 0xeb
    x"00000000", -- 236, 0xec
    x"00000000", -- 237, 0xed
    x"00000000", -- 238, 0xee
    x"00000000", -- 239, 0xef
    x"00000000", -- 240, 0xf0
    x"00000000", -- 241, 0xf1
    x"00000000", -- 242, 0xf2
    x"00000000", -- 243, 0xf3
    x"00000000", -- 244, 0xf4
    x"00000000", -- 245, 0xf5
    x"00000000", -- 246, 0xf6
    x"00000000", -- 247, 0xf7
    x"00000000", -- 248, 0xf8
    x"00000000", -- 249, 0xf9
    x"00000000", -- 250, 0xfa
    x"00000000", -- 251, 0xfb
    x"00000000", -- 252, 0xfc
    x"00000000", -- 253, 0xfd
    x"00000000", -- 254, 0xfe
    x"00000000" -- 255, 0xff
    );
    signal sarr256lv32_hash_table_memory_0 : hash_table_memory_t := (-- LSW
    x"00000000", -- 0, 0x00
    x"00000000", -- 1, 0x01
    x"00000000", -- 2, 0x02
    x"00000000", -- 3, 0x03
    x"00000000", -- 4, 0x04
    x"00000000", -- 5, 0x05
    x"00000000", -- 6, 0x06
    x"00000000", -- 7, 0x07
    x"00000000", -- 8, 0x08
    x"00000000", -- 9, 0x09
    x"00000000", -- 10, 0x0a
    x"00000000", -- 11, 0x0b
    x"00000000", -- 12, 0x0c
    x"00000000", -- 13, 0x0d
    x"00000000", -- 14, 0x0e
    x"00000000", -- 15, 0x0f
    x"00000000", -- 16, 0x10
    x"00000000", -- 17, 0x11
    x"00000000", -- 18, 0x12
    x"00000000", -- 19, 0x13
    x"00000000", -- 20, 0x14
    x"00000000", -- 21, 0x15
    x"00000000", -- 22, 0x16
    x"00000000", -- 23, 0x17
    x"00000000", -- 24, 0x18
    x"00000000", -- 25, 0x19
    x"00000000", -- 26, 0x1a
    x"00000000", -- 27, 0x1b
    x"00000000", -- 28, 0x1c
    x"00000000", -- 29, 0x1d
    x"00000000", -- 30, 0x1e
    x"00000000", -- 31, 0x1f
    x"00000000", -- 32, 0x20
    x"00000000", -- 33, 0x21
    x"00000000", -- 34, 0x22
    x"00000000", -- 35, 0x23
    x"00000000", -- 36, 0x24
    x"00000000", -- 37, 0x25
    x"00000000", -- 38, 0x26
    x"00000000", -- 39, 0x27
    x"00000000", -- 40, 0x28
    x"00000000", -- 41, 0x29
    x"00000000", -- 42, 0x2a
    x"00000000", -- 43, 0x2b
    x"00000000", -- 44, 0x2c
    x"00000000", -- 45, 0x2d
    x"00000000", -- 46, 0x2e
    x"00000000", -- 47, 0x2f
    x"00000000", -- 48, 0x30
    x"00000000", -- 49, 0x31
    x"00000000", -- 50, 0x32
    x"00000000", -- 51, 0x33
    x"00000000", -- 52, 0x34
    x"00000000", -- 53, 0x35
    x"00000000", -- 54, 0x36
    x"00000000", -- 55, 0x37
    x"00000000", -- 56, 0x38
    x"00000000", -- 57, 0x39
    x"00000000", -- 58, 0x3a
    x"00000000", -- 59, 0x3b
    x"00000000", -- 60, 0x3c
    x"00000000", -- 61, 0x3d
    x"00000000", -- 62, 0x3e
    x"00000000", -- 63, 0x3f
    x"00000000", -- 64, 0x40
    x"00000000", -- 65, 0x41
    x"00000000", -- 66, 0x42
    x"00000000", -- 67, 0x43
    x"00000000", -- 68, 0x44
    x"00000000", -- 69, 0x45
    x"00000000", -- 70, 0x46
    x"00000000", -- 71, 0x47
    x"00000000", -- 72, 0x48
    x"00000000", -- 73, 0x49
    x"00000000", -- 74, 0x4a
    x"00000000", -- 75, 0x4b
    x"00000000", -- 76, 0x4c
    x"00000000", -- 77, 0x4d
    x"00000000", -- 78, 0x4e
    x"00000000", -- 79, 0x4f
    x"00000000", -- 80, 0x50
    x"00000000", -- 81, 0x51
    x"00000000", -- 82, 0x52
    x"00000000", -- 83, 0x53
    x"00000000", -- 84, 0x54
    x"00000000", -- 85, 0x55
    x"00000000", -- 86, 0x56
    x"00000000", -- 87, 0x57
    x"00000000", -- 88, 0x58
    x"00000000", -- 89, 0x59
    x"00000000", -- 90, 0x5a
    x"00000000", -- 91, 0x5b
    x"00000000", -- 92, 0x5c
    x"00000000", -- 93, 0x5d
    x"00000000", -- 94, 0x5e
    x"00000000", -- 95, 0x5f
    x"00000000", -- 96, 0x60
    x"00000000", -- 97, 0x61
    x"00000000", -- 98, 0x62
    x"00000000", -- 99, 0x63
    x"00000000", -- 100, 0x64
    x"00000000", -- 101, 0x65
    x"00000000", -- 102, 0x66
    x"00000000", -- 103, 0x67
    x"00000000", -- 104, 0x68
    x"00000000", -- 105, 0x69
    x"00000000", -- 106, 0x6a
    x"00000000", -- 107, 0x6b
    x"00000000", -- 108, 0x6c
    x"00000000", -- 109, 0x6d
    x"00000000", -- 110, 0x6e
    x"00000000", -- 111, 0x6f
    x"00000000", -- 112, 0x70
    x"00000000", -- 113, 0x71
    x"00000000", -- 114, 0x72
    x"00000000", -- 115, 0x73
    x"00000000", -- 116, 0x74
    x"00000000", -- 117, 0x75
    x"00000000", -- 118, 0x76
    x"00000000", -- 119, 0x77
    x"00000000", -- 120, 0x78
    x"00000000", -- 121, 0x79
    x"00000000", -- 122, 0x7a
    x"00000000", -- 123, 0x7b
    x"00000000", -- 124, 0x7c
    x"00000000", -- 125, 0x7d
    x"00000000", -- 126, 0x7e
    x"00000000", -- 127, 0x7f
    x"00000000", -- 128, 0x80
    x"00000000", -- 129, 0x81
    x"00000000", -- 130, 0x82
    x"00000000", -- 131, 0x83
    x"00000000", -- 132, 0x84
    x"00000000", -- 133, 0x85
    x"00000000", -- 134, 0x86
    x"00000000", -- 135, 0x87
    x"00000000", -- 136, 0x88
    x"00000000", -- 137, 0x89
    x"00000000", -- 138, 0x8a
    x"00000000", -- 139, 0x8b
    x"00000000", -- 140, 0x8c
    x"00000000", -- 141, 0x8d
    x"00000000", -- 142, 0x8e
    x"00000000", -- 143, 0x8f
    x"00000000", -- 144, 0x90
    x"00000000", -- 145, 0x91
    x"00000000", -- 146, 0x92
    x"00000000", -- 147, 0x93
    x"00000000", -- 148, 0x94
    x"00000000", -- 149, 0x95
    x"00000000", -- 150, 0x96
    x"00000000", -- 151, 0x97
    x"00000000", -- 152, 0x98
    x"00000000", -- 153, 0x99
    x"00000000", -- 154, 0x9a
    x"00000000", -- 155, 0x9b
    x"00000000", -- 156, 0x9c
    x"00000000", -- 157, 0x9d
    x"00000000", -- 158, 0x9e
    x"00000000", -- 159, 0x9f
    x"00000000", -- 160, 0xa0
    x"00000000", -- 161, 0xa1
    x"00000000", -- 162, 0xa2
    x"00000000", -- 163, 0xa3
    x"00000000", -- 164, 0xa4
    x"00000000", -- 165, 0xa5
    x"00000000", -- 166, 0xa6
    x"00000000", -- 167, 0xa7
    x"00000000", -- 168, 0xa8
    x"00000000", -- 169, 0xa9
    x"00000000", -- 170, 0xaa
    x"00000000", -- 171, 0xab
    x"00000000", -- 172, 0xac
    x"00000000", -- 173, 0xad
    x"00000000", -- 174, 0xae
    x"00000000", -- 175, 0xaf
    x"00000000", -- 176, 0xb0
    x"00000000", -- 177, 0xb1
    x"00000000", -- 178, 0xb2
    x"00000000", -- 179, 0xb3
    x"00000000", -- 180, 0xb4
    x"00000000", -- 181, 0xb5
    x"00000000", -- 182, 0xb6
    x"00000000", -- 183, 0xb7
    x"00000000", -- 184, 0xb8
    x"00000000", -- 185, 0xb9
    x"00000000", -- 186, 0xba
    x"00000000", -- 187, 0xbb
    x"00000000", -- 188, 0xbc
    x"00000000", -- 189, 0xbd
    x"00000000", -- 190, 0xbe
    x"00000000", -- 191, 0xbf
    x"00000000", -- 192, 0xc0
    x"00000000", -- 193, 0xc1
    x"00000000", -- 194, 0xc2
    x"00000000", -- 195, 0xc3
    x"00000000", -- 196, 0xc4
    x"00000000", -- 197, 0xc5
    x"00000000", -- 198, 0xc6
    x"67000000", -- 199, 0xc7
    x"00000000", -- 200, 0xc8
    x"00000000", -- 201, 0xc9
    x"00000000", -- 202, 0xca
    x"00000000", -- 203, 0xcb
    x"00000000", -- 204, 0xcc
    x"00000000", -- 205, 0xcd
    x"00000000", -- 206, 0xce
    x"00000000", -- 207, 0xcf
    x"00000000", -- 208, 0xd0
    x"00000000", -- 209, 0xd1
    x"00000000", -- 210, 0xd2
    x"00000000", -- 211, 0xd3
    x"00000000", -- 212, 0xd4
    x"00000000", -- 213, 0xd5
    x"00000000", -- 214, 0xd6
    x"00000000", -- 215, 0xd7
    x"00000000", -- 216, 0xd8
    x"00000000", -- 217, 0xd9
    x"00000000", -- 218, 0xda
    x"00000000", -- 219, 0xdb
    x"00000000", -- 220, 0xdc
    x"00000000", -- 221, 0xdd
    x"00000000", -- 222, 0xde
    x"00000000", -- 223, 0xdf
    x"00000000", -- 224, 0xe0
    x"00000000", -- 225, 0xe1
    x"FF000000", -- 226, 0xe2
    x"00000000", -- 227, 0xe3
    x"00000000", -- 228, 0xe4
    x"00000000", -- 229, 0xe5
    x"00000000", -- 230, 0xe6
    x"00000000", -- 231, 0xe7
    x"00000000", -- 232, 0xe8
    x"00000000", -- 233, 0xe9
    x"00000000", -- 234, 0xea
    x"00000000", -- 235, 0xeb
    x"00000000", -- 236, 0xec
    x"00000000", -- 237, 0xed
    x"00000000", -- 238, 0xee
    x"00000000", -- 239, 0xef
    x"00000000", -- 240, 0xf0
    x"00000000", -- 241, 0xf1
    x"00000000", -- 242, 0xf2
    x"00000000", -- 243, 0xf3
    x"00000000", -- 244, 0xf4
    x"00000000", -- 245, 0xf5
    x"00000000", -- 246, 0xf6
    x"00000000", -- 247, 0xf7
    x"00000000", -- 248, 0xf8
    x"00000000", -- 249, 0xf9
    x"00000000", -- 250, 0xfa
    x"00000000", -- 251, 0xfb
    x"00000000", -- 252, 0xfc
    x"00000000", -- 253, 0xfd
    x"00000000", -- 254, 0xfe
    x"00000000" -- 255, 0xff
    );
    signal slv32_hash_table_rd_data_3 : std_logic_vector(ACL_HASH_TABLE_M9K_LENGTH - 1 downto 0) := (others => '0');
    signal slv32_hash_table_rd_data_2 : std_logic_vector(ACL_HASH_TABLE_M9K_LENGTH - 1 downto 0) := (others => '0');
    signal slv32_hash_table_rd_data_1 : std_logic_vector(ACL_HASH_TABLE_M9K_LENGTH - 1 downto 0) := (others => '0');
    signal slv32_hash_table_rd_data_0 : std_logic_vector(ACL_HASH_TABLE_M9K_LENGTH - 1 downto 0) := (others => '0');

    -- signal slv32_hash_table_wr_data_3 : std_logic_vector(ACL_HASH_TABLE_M9K_LENGTH - 1 downto 0) := (others => '0');
    -- signal slv32_hash_table_wr_data_2 : std_logic_vector(ACL_HASH_TABLE_M9K_LENGTH - 1 downto 0) := (others => '0');
    -- signal slv32_hash_table_wr_data_1 : std_logic_vector(ACL_HASH_TABLE_M9K_LENGTH - 1 downto 0) := (others => '0');
    -- signal slv32_hash_table_wr_data_0 : std_logic_vector(ACL_HASH_TABLE_M9K_LENGTH - 1 downto 0) := (others => '0');
begin
    --    slv32_hash_table_wr_data_3 <= pilv128_hash_wr_value(ACL_HASH_TABLE_M9K_LENGTH * 4 - 1 downto ACL_HASH_TABLE_M9K_LENGTH * 3);
    --    slv32_hash_table_wr_data_2 <= pilv128_hash_wr_value(ACL_HASH_TABLE_M9K_LENGTH * 3 - 1 downto ACL_HASH_TABLE_M9K_LENGTH * 2);
    --    slv32_hash_table_wr_data_1 <= pilv128_hash_wr_value(ACL_HASH_TABLE_M9K_LENGTH * 2 - 1 downto ACL_HASH_TABLE_M9K_LENGTH * 1);
    --    slv32_hash_table_wr_data_0 <= pilv128_hash_wr_value(ACL_HASH_TABLE_M9K_LENGTH * 1 - 1 downto 0);
    --
    polv128_hash_rd_value <= slv32_hash_table_rd_data_3 &
        slv32_hash_table_rd_data_2 &
        slv32_hash_table_rd_data_1 &
        slv32_hash_table_rd_data_0;

    process (pil_clk)
    begin
        if rising_edge(pil_clk) then
            --    if (pil_hash_wr_en = '1') then
            --
            --        sarr256lv32_hash_table_memory_3(to_integer(unsigned(pilv8_hash_table_wr_addr))) <= slv32_hash_table_wr_data_3;
            --        sarr256lv32_hash_table_memory_2(to_integer(unsigned(pilv8_hash_table_wr_addr))) <= slv32_hash_table_wr_data_2;
            --        sarr256lv32_hash_table_memory_1(to_integer(unsigned(pilv8_hash_table_wr_addr))) <= slv32_hash_table_wr_data_1;
            --        sarr256lv32_hash_table_memory_0(to_integer(unsigned(pilv8_hash_table_wr_addr))) <= slv32_hash_table_wr_data_0;
            --
            --    end if;
            if (pil_hash_rd_en = '1') then
                slv32_hash_table_rd_data_3 <= sarr256lv32_hash_table_memory_3(to_integer(unsigned(pilv8_hash_table_rd_addr)));
                slv32_hash_table_rd_data_2 <= sarr256lv32_hash_table_memory_2(to_integer(unsigned(pilv8_hash_table_rd_addr)));
                slv32_hash_table_rd_data_1 <= sarr256lv32_hash_table_memory_1(to_integer(unsigned(pilv8_hash_table_rd_addr)));
                slv32_hash_table_rd_data_0 <= sarr256lv32_hash_table_memory_0(to_integer(unsigned(pilv8_hash_table_rd_addr)));
            else

            end if;
        end if;
    end process;
end architecture;